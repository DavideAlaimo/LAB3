library ieee;
use ieee.std_logic_1164.all;

ENTITY ZeroGenerating IS
PORT (OUT_REG1,OUT_REG2,BYPASS_ALU,BYPASS_WB : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      OPCODE_1 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
      SEL_MUX_ALU_SRC1, SEL_MUX_ALU_SRC2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      FLAG_FORWARDING_A, FLAG_FORWARDING_B : IN STD_LOGIC;
      ZERO_GENERATED : OUT STD_LOGIC
      );
END ENTITY;

ARCHITECTURE BEH OF ZeroGenerating IS

COMPONENT COMPARE IS
PORT (IN1, IN2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      OUT_COMPARE : OUT STD_LOGIC);
END COMPONENT;

SIGNAL COMP_REG1_REG2, COMP_REG1_BYPASS_ALU, COMP_REG1_BYPASS_WB,
        COMP_REG2_BYPASS_ALU, COMP_REG2_BYPASS_WB :STD_LOGIC;

BEGIN

COMPARE_REG1_REG2 : COMPARE PORT MAP(OUT_REG1,OUT_REG2,COMP_REG1_REG2);
COMPARE_REG1_BYPASS_ALU : COMPARE PORT MAP(OUT_REG1,BYPASS_ALU,COMP_REG1_BYPASS_ALU);
COMPARE_REG1_BYPASS_WB : COMPARE PORT MAP(OUT_REG1,BYPASS_WB,COMP_REG1_BYPASS_WB);
COMPARE_REG2_BYPASS_ALU : COMPARE PORT MAP(OUT_REG2,BYPASS_ALU,COMP_REG2_BYPASS_ALU);
COMPARE_REG2_BYPASS_WB : COMPARE PORT MAP(OUT_REG2,BYPASS_WB,COMP_REG2_BYPASS_WB);

PROCESS(OPCODE_1,SEL_MUX_ALU_SRC1,SEL_MUX_ALU_SRC2,FLAG_FORWARDING_A,FLAG_FORWARDING_B,
	COMP_REG1_REG2,COMP_REG1_BYPASS_ALU,COMP_REG1_BYPASS_WB,COMP_REG2_BYPASS_ALU,COMP_REG2_BYPASS_WB) 
VARIABLE CASE_SELECTOR: STD_LOGIC_VECTOR(14 DOWNTO 0);
VARIABLE OUT_COMPARE:STD_LOGIC;
BEGIN
CASE_SELECTOR := OPCODE_1 & SEL_MUX_ALU_SRC1 & SEL_MUX_ALU_SRC2 & FLAG_FORWARDING_A & FLAG_FORWARDING_B;
CASE (CASE_SELECTOR) IS 

--OPCODE_1="1100011"; SEL_MUX_ALU_SRC1="000"; SEL_MUX_ALU_SRC2="000"; FLAG_FORWARDING_A='0'; FLAG_FORWARDING_B='0'
WHEN ("110001100000000") => ZERO_GENERATED<=COMP_REG1_REG2;

--OPCODE_1="1100011"; SEL_MUX_ALU_SRC1="000"; SEL_MUX_ALU_SRC2="011"; FLAG_FORWARDING_A='0'; FLAG_FORWARDING_B='1'
WHEN ("110001100001101") => ZERO_GENERATED<=COMP_REG1_BYPASS_ALU;

--OPCODE_1="1100011"; SEL_MUX_ALU_SRC1="000"; SEL_MUX_ALU_SRC2="100"; FLAG_FORWARDING_A='0'; FLAG_FORWARDING_B='1'
WHEN ("110001100010001") => ZERO_GENERATED<=COMP_REG1_BYPASS_WB;

--OPCODE_1="1100011"; SEL_MUX_ALU_SRC1="011"; SEL_MUX_ALU_SRC2="000"; FLAG_FORWARDING_A='1'; FLAG_FORWARDING_B='0'
WHEN ("110001101100010") => ZERO_GENERATED<=COMP_REG2_BYPASS_ALU;

--OPCODE_1="1100011"; SEL_MUX_ALU_SRC1="100"; SEL_MUX_ALU_SRC2="000"; FLAG_FORWARDING_A='1'; FLAG_FORWARDING_B='0'
WHEN ("110001110000010") => ZERO_GENERATED<=COMP_REG2_BYPASS_WB;

WHEN OTHERS => ZERO_GENERATED<='0';

END CASE;

END PROCESS;
END ARCHITECTURE;