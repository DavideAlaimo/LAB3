library ieee;
use ieee.std_logic_1164.all;

ENTITY Reg IS
PORT(DATA_IN : IN STD_LOGIC;
     CLK, RST: IN STD_LOGIC;
     DATA_OUT : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEH OF Reg IS
BEGIN
PROCESS(CLK, RST)
BEGIN
IF(RST='1') THEN DATA_OUT<='0'; 
ELSIF(CLK'event  and  CLK='1') THEN  DATA_OUT<=DATA_IN;
END IF;
END PROCESS;
END ARCHITECTURE;