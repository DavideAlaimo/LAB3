library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;



ENTITY ControlHazardUnit2 IS
PORT(OPCODE_1: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
	ZERO_ALU,CLK,RST: IN STD_LOGIC;
	SEL_MUX_PC,SEL_MUX_INSTR: OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEH OF ControlHazardUnit2 IS

--TYPE STATE IS (IDLE,S1);
--SIGNAL PSTATE,NSTATE : STATE;
SIGNAL STATE : STD_LOGIC; --0 IDLE 1 S1
SIGNAL PSTATE,NSTATE : STD_LOGIC;
SIGNAL BEQ_CONDITION : STD_LOGIC;
SIGNAL MUX_PC_ASM,MUX_PC_DT, MUX_INSTR_ASM, MUX_INSTR_DT : STD_LOGIC;
--SIGNAL MUX_PC_RST,MUX_INSTR_RST:STD_LOGIC;

COMPONENT Reg IS
PORT(DATA_IN : IN STD_LOGIC;
     CLK, RST: IN STD_LOGIC;
     DATA_OUT : OUT STD_LOGIC);
END COMPONENT;

BEGIN
BEQ_CONDITION <= '1' WHEN OPCODE_1="1100011" AND ZERO_ALU='1' ELSE '0';
--MUX_PC_ASM<='0';MUX_PC_DT<='0'; MUX_INSTR_ASM<='0'; MUX_INSTR_DT<='0';
--MUX_PC_RST<='0';MUX_INSTR_RST<='0';


--    PROCESS(CLK,RST)
--      BEGIN
--        IF(RST='1') THEN PSTATE<='0';--MUX_PC_DT<='0'; MUX_INSTR_DT<='0';
--        ELSIF (CLK'EVENT AND CLK='1') THEN PSTATE<=NSTATE;
--        END IF;
--    END PROCESS;

PSTATE_REGISTER : Reg PORT MAP(NSTATE,CLK,RST,PSTATE);

PROCESS(PSTATE,BEQ_CONDITION)

BEGIN
CASE (PSTATE) IS
	WHEN '0' =>   IF(BEQ_CONDITION='1') THEN NSTATE<='1'; 
			ELSIF(BEQ_CONDITION='0') THEN  NSTATE<='0'; 
			END IF;
	WHEN '1' => NSTATE<='0'; 
	WHEN OTHERS => NSTATE<='1'; 
END CASE;
END PROCESS;

MUX_PC_DT <='1' WHEN BEQ_CONDITION='1' ELSE '0';
MUX_INSTR_DT <='1' WHEN BEQ_CONDITION='1' ELSE '0';

SEL_MUX_PC <= MUX_PC_DT OR MUX_PC_ASM;-- OR MUX_PC_RST;
SEL_MUX_INSTR <= MUX_INSTR_DT OR MUX_INSTR_ASM;--OR MUX_INSTR_RST;

PROCESS(PSTATE) 
BEGIN
CASE(PSTATE) IS
	WHEN '0' => MUX_PC_ASM<='0'; MUX_INSTR_ASM<='0'; 
	WHEN '1' =>   MUX_PC_ASM<='0'; MUX_INSTR_ASM<='0';
	WHEN OTHERS => MUX_PC_ASM<='0'; MUX_INSTR_ASM<='0';
END CASE;
END PROCESS;

END ARCHITECTURE;