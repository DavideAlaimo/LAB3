library ieee;
use ieee.std_logic_1164.all;

ENTITY COMPARE IS
PORT (IN1, IN2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      OUT_COMPARE : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEH OF COMPARE IS

BEGIN
PROCESS(IN1,IN2) 
BEGIN
IF (IN1=IN2) THEN OUT_COMPARE <= '1';
ELSE OUT_COMPARE <= '0';
END IF;
END PROCESS;

END ARCHITECTURE;
