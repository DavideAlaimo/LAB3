library ieee;
use ieee.std_logic_1164.all;

ENTITY MUX_5TO1 IS
PORT(IN1,IN2,IN3,IN4,IN5 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     SELECTOR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
     OUT_MUX_5TO1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEH OF MUX_5TO1 IS
BEGIN
PROCESS(SELECTOR,IN1,IN2,IN3,IN4,IN5)
BEGIN
IF(SELECTOR="000") THEN OUT_MUX_5TO1 <= IN1;
ELSIF(SELECTOR="001") THEN OUT_MUX_5TO1 <= IN2;
ELSIF(SELECTOR="010") THEN OUT_MUX_5TO1 <= IN3;
ELSIF(SELECTOR="011") THEN OUT_MUX_5TO1 <= IN4; -- FORWARD A EX_MEM
ELSIF(SELECTOR="100") THEN OUT_MUX_5TO1 <= IN5; -- FORWARD B MEM_WB
ELSE OUT_MUX_5TO1 <= (OTHERS=>'U');
END IF;
END PROCESS;
END ARCHITECTURE;
