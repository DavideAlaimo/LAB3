library ieee;
use ieee.std_logic_1164.all;

ENTITY MUX_2TO1 IS
GENERIC (N : INTEGER );
PORT(IN1,IN2 : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
     SELECTOR : IN STD_LOGIC;
     OUT_MUX_2TO1 : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEH OF MUX_2TO1 IS
BEGIN
PROCESS(SELECTOR,IN1,IN2)
BEGIN
IF(SELECTOR='0') THEN OUT_MUX_2TO1 <= IN1;
ELSIF(SELECTOR='1') THEN OUT_MUX_2TO1 <= IN2;
ELSE OUT_MUX_2TO1 <= (OTHERS=>'U');
END IF;
END PROCESS;
END ARCHITECTURE;