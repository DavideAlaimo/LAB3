library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all; 

ENTITY RISC_V IS
PORT(INSTRUCTION : IN STD_LOGIC_VECTOR(31 DOWNTO 0); --DATA OUTPUT MEMORY INSTRUCTION
     DATA_OUT_MEM_DATA : IN STD_LOGIC_VECTOR(63 DOWNTO 0); -- DATA OUTPUT MEMORY DATA
     CLK, RST : IN STD_LOGIC;
     ADDRESS_MEM_INSTR, ADDRESS_MEM_DATA : OUT STD_LOGIC_VECTOR(63 DOWNTO 0); --ADDRESSES DATA AND INSTRUCTION MEMORY
     DATA_TOWRITE_MEM_DATA : OUT STD_LOGIC_VECTOR(63 DOWNTO 0); --DATA TO WRITE IN MEMORY DATA
     READ_MEM_DATA, WRITE_MEM_DATA,EN_ISTR_MEM : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE BEH OF RISC_V IS

--ADDER TO COMPUTE NEXT ADDRESS SEQUENTIAL OR JUMP
COMPONENT Adder IS   
GENERIC (N : INTEGER :=64);
PORT(IN1, IN2 : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
     RST : IN STD_LOGIC;
     OUT_SUM : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;

COMPONENT ALU IS
PORT(IN1, IN2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     OP: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
     Zero : OUT STD_LOGIC;
     OUT_ALU : BUFFER STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT AluControl IS
PORT(ALUop : IN STD_LOGIC;
     INSTR30 : IN STD_LOGIC;
     FUNCT3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
     ALUoperation : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END COMPONENT;

COMPONENT CONTROL IS
PORT(OPCODE : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
     RD:IN STD_LOGIC_VECTOR(4 DOWNTO 0);
     Branch, MemRead, MemToReg, ALUop, MemWrite, RegWrite, MuxToBranch : OUT STD_LOGIC;
     ALUsrc1, ALUsrc2 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
     EnFunctUnit : OUT STD_LOGIC);
END COMPONENT;

COMPONENT ImmediateGenerator IS
PORT (Instruction : IN STD_LOGIC_VECTOR(31 downto 0);
      Instruction_64 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT MUX_2TO1 IS
GENERIC (N : INTEGER );
PORT(IN1,IN2 : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
     SELECTOR : IN STD_LOGIC;
     OUT_MUX_2TO1 : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));
END COMPONENT;

COMPONENT MUX_5TO1 IS
PORT(IN1,IN2,IN3,IN4,IN5 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     SELECTOR : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
     OUT_MUX_5TO1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT ForwardingUnit IS
PORT(RS1,RS2,RD_EX_MEM,RD_MEM_WB : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
     RegWrite_EX_MEM, RegWrite_MEM_WB : IN STD_LOGIC; 
     ForwardA, ForwardB : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
     PriorityA, PriorityB : OUT STD_LOGIC);
END COMPONENT;

COMPONENT  HazardDetectionUnit IS
PORT(	RS1,RS2,RD,WriteReg : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	RegWrite,MemRead,Foreward_on,CLK: IN STD_LOGIC;
	EN_PC, EN_IF_ID,EN_ID_EX: OUT STD_LOGIC;
	MUX_BUBBLE: OUT STD_LOGIC);
END COMPONENT;

COMPONENT ZeroGenerating IS
PORT (OUT_REG1,OUT_REG2,BYPASS_ALU,BYPASS_WB : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      OPCODE_1 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
      SEL_MUX_ALU_SRC1, SEL_MUX_ALU_SRC2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      FLAG_FORWARDING_A, FLAG_FORWARDING_B : IN STD_LOGIC;
      ZERO_GENERATED : OUT STD_LOGIC
      );
END COMPONENT;

COMPONENT FunctionUnit IS
PORT(EN_FUNCT : IN STD_LOGIC;
     DATA_IN : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     DATA_OUT : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT Register_N IS
PORT(DATA_IN : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     CLK, RST, EN : IN STD_LOGIC;
     DATA_OUT : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT PC_Register IS

PORT(DATA_IN : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
     CLK, RST, EN : IN STD_LOGIC;
     DATA_OUT : OUT STD_LOGIC_VECTOR(63 DOWNTO 0));
END COMPONENT;

COMPONENT RegistersFile IS
PORT(ReadReg1, ReadReg2, WriteReg  : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    WriteData : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    CLK, RegWrite, RST : IN STD_LOGIC;
    ReadData1, ReadData2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
     );
END COMPONENT;

COMPONENT ControlHazardUnit IS
	PORT(OPCODE,OPCODE_1: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
	     ZERO_ALU,CLK,RST: IN STD_LOGIC;		
	SEL_MUX_PC,SEL_MUX_INSTR: OUT STD_LOGIC);
END COMPONENT;




---------------------------------------------------SIGNALS------------------------------------------------------------------
---------------------- SIGNALS CONTROL UNIT
SIGNAL SIGNALS_CONTROL, NEW_SIGNALS_CONTROL : STD_LOGIC_VECTOR(13 DOWNTO 0);
SIGNAL BRANCH, MEM_READ, MEM_WRITE, MEM_TO_REG, ALUop, REG_WRITE, MUX_TO_BRANCH : STD_LOGIC;
SIGNAL ALU_src1, ALU_src2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL BRANCH0, MEM_READ0, MEM_WRITE0, MEM_TO_REG0, ALUop0, REG_WRITE0, MUX_TO_BRANCH0 : STD_LOGIC;
SIGNAL ALU_src10, ALU_src20 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL EN_PC, EN_IF_ID, MUX_SEL_BUBBLE : STD_LOGIC;
SIGNAL EN_FUNCT0, EN_FUNCT : STD_LOGIC;
--FIRST LEVEL PIPE
SIGNAL BRANCH1, MEM_READ1, MEM_WRITE1, MEM_TO_REG1, ALUop1, REG_WRITE1, MUX_TO_BRANCH1 : STD_LOGIC;
SIGNAL ALU_src11, ALU_src21  : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL EN_FUNCT1 : STD_LOGIC;
--SECOND LEVEL PIPE
SIGNAL BRANCH2, MEM_TO_REG2, REG_WRITE2, MUX_TO_BRANCH2 : STD_LOGIC;
--THIRD LEVEL PIPE
SIGNAL MEM_TO_REG3, REG_WRITE3: STD_LOGIC;


---------------------DATAPATH SIGNALS
SIGNAL OUT_PC : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_ADD_SEQUENTIAL : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_ADD_BRANCH : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_REG_FILE1, OUT_REG_FILE2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_IMM_GEN : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_MUX_SRC1, OUT_MUX_SRC2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_ALU_CONTROL : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL OUT_ZERO_ALU : STD_LOGIC; SIGNAL OUT_RESULT_ALU : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_MUX_BRANCH : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL OUT_MUX_MEM_TO_REG : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_MUX_SEQ_BRANCH : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_REG0, OUT_REG4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_INSTR_FUNCT : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL OUT_IMM_GEN_1_SHIFTED : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL SELECTOR_MUX_BRANCH_SEQ : STD_LOGIC;
SIGNAL ADD_REG_WRITE : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL OUT_COMPARATOR : STD_LOGIC;
SIGNAL OUT_FUNCT : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_MUX_FUNCT_ALU : STD_LOGIC_VECTOR(63 DOWNTO 0);

-------------------SIGNAL HAZARD/COUNTER

SIGNAL CNT: UNSIGNED(1 DOWNTO 0);
SIGNAL EN_CNT, EN_ID_EX: STD_LOGIC;
SIGNAL RST_CNT_HZ: STD_LOGIC;
SIGNAL RST_CNT :STD_LOGIC;
SIGNAL TC: STD_LOGIC;
SIGNAL MUX_PC:STD_LOGIC;
SIGNAL OUT_MUX_PC:STD_LOGIC_VECTOR(63 DOWNTO 0);



-------------------DATAPATH PIPE SIGNALS

SIGNAL RS1,RS1_1,RS2,RS2_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL RD, RD_1, RD_2_EX_MEM, RD_3_MEM_WB : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL FORWARD_A, FORWARD_B : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL FA_FLAG, FB_FLAG : STD_LOGIC; 
SIGNAL NEW_MUX_SRC1_SEL, NEW_MUX_SRC2_SEL : STD_LOGIC_VECTOR(2 DOWNTO 0);


--FIRST PIPE LEVEL : OUT ADDER SEQUENTIAL, OUT PC, OUT INSTRUCTION

SIGNAL OUT_PC_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL INSTRUCTION_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);


--SECOND PIPE LEVEL : READ DATA 1, READ DATA 2, OUT IMM GEN, OUT INSTR FUNCT 3, OUT ADDER SEQUENTIAL PIPE 1, OUT PC PIPE 1, OUT REG '0', OUT REG 4

SIGNAL MUX_INSTR: STD_LOGIC;
SIGNAL OPCODE_1: STD_lOGIC_VECTOR(6 DOWNTO 0);
SIGNAL OUT_PC_2, OUT_REG0_1, OUT_REG4_1,  OUT_REG_FILE1_1, OUT_REG_FILE2_1, OUT_IMM_GEN_1: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_INSTR_FUNCT_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL ADD_REG_WRITE_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL Forward_on:std_logic;


--THIRD LEVEL PIPE : OUT ADDER SEQUENTIAL PIPE 2, OUT ADDER BRANCH, OUT ALU ZERO, OUT ALU RESULT, READ DATA 2, SIGNAL OUT_PC_3

SIGNAL OUT_ADD_BRANCH_1, OUT_RESULT_ALU_1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_ZERO_ALU_1 : STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL ADD_REG_WRITE_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);


--FOURTH LEVEL PIPE : OUT MEMORY DATA, OUT ALU RESULT PIPE 1

SIGNAL DATA_OUT_MEM_DATA_1: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL OUT_RESULT_ALU_2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL ADD_REG_WRITE_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);


BEGIN



PC : PC_Register PORT MAP (OUT_MUX_SEQ_BRANCH, CLK, RST,EN_PC, OUT_PC);

ZERO_GENERATING_COMPONENT : ZeroGenerating PORT MAP(OUT_REG_FILE1_1,OUT_REG_FILE2_1,OUT_RESULT_ALU_1,OUT_MUX_MEM_TO_REG,
OPCODE_1,NEW_MUX_SRC1_SEL,NEW_MUX_SRC2_SEL,FA_FLAG,FB_FLAG,OUT_COMPARATOR);

MuxPC : MUX_2TO1 GENERIC MAP(64) PORT MAP(OUT_PC, x"0000000000400054", MUX_PC, OUT_MUX_PC);

ADDRESS_MEM_INSTR<=OUT_MUX_PC;

ADDER_SEQUENTIAL : Adder PORT MAP (OUT_MUX_PC, x"0000000000000004", RST, OUT_ADD_SEQUENTIAL);

ADDER_JUMP : Adder PORT MAP (OUT_PC_2, OUT_IMM_GEN_1_SHIFTED, RST, OUT_ADD_BRANCH);

Registers_File : RegistersFile PORT MAP (INSTRUCTION_1(19 DOWNTO 15), INSTRUCTION_1(24 DOWNTO 20), ADD_REG_WRITE_2, OUT_MUX_MEM_TO_REG, CLK, REG_WRITE3, RST, OUT_REG_FILE1, OUT_REG_FILE2);

IMMEDIATE_GENERATOR : ImmediateGenerator PORT MAP (INSTRUCTION_1, OUT_IMM_GEN);

MuxINSTR : MUX_2TO1 GENERIC MAP(32) PORT MAP(INSTRUCTION, x"00000013", MUX_INSTR, INSTRUCTION_1);

ControlHZ: ControlHazardUnit PORT MAP(INSTRUCTION_1(6 DOWNTO 0),OPCODE_1,OUT_COMPARATOR,CLK,RST,MUX_PC,MUX_INSTR);

--LEFT SHIFT OUT_IMM_GEN_1
PROCESS(OUT_IMM_GEN_1)

VARIABLE IMM_SIGNED : SIGNED (63 DOWNTO 0);
VARIABLE OUT_SHIFT : SIGNED(63 DOWNTO 0);

BEGIN

IMM_SIGNED := SIGNED(OUT_IMM_GEN_1);
OUT_SHIFT := SHIFT_LEFT(IMM_SIGNED,1);
OUT_IMM_GEN_1_SHIFTED <= STD_LOGIC_VECTOR(OUT_SHIFT);

END PROCESS;

ALU_CONTROL : AluControl PORT MAP(ALUop1, INSTRUCTION_1(30), OUT_INSTR_FUNCT_1, OUT_ALU_CONTROL);

ALU_COMPONENT : ALU PORT MAP(OUT_MUX_SRC1, OUT_MUX_SRC2, OUT_ALU_CONTROL, OUT_ZERO_ALU, OUT_RESULT_ALU);

SPECIAL_FUNCTION_UNIT : FunctionUnit PORT MAP(EN_FUNCT1,OUT_MUX_SRC1,OUT_FUNCT);

MUX_FUNCT_OR_ALU : MUX_2TO1 GENERIC MAP(64) PORT MAP(OUT_RESULT_ALU,OUT_FUNCT,EN_FUNCT1,OUT_MUX_FUNCT_ALU);

CONTROL_UNIT : CONTROL PORT MAP (INSTRUCTION_1(6 DOWNTO 0),INSTRUCTION_1(11 DOWNTO 7), BRANCH0, MEM_READ0, MEM_TO_REG0, ALUop0, MEM_WRITE0, REG_WRITE0, MUX_TO_BRANCH0, ALU_src10, ALU_src20,EN_FUNCT0);

SIGNALS_CONTROL <= EN_FUNCT0&BRANCH0&MEM_READ0&MEM_TO_REG0&ALUop0&MEM_WRITE0&REG_WRITE0&MUX_TO_BRANCH0&ALU_src10&ALU_src20;

MUX_ALU_SRC1 : MUX_5TO1 PORT MAP(OUT_REG_FILE1_1, OUT_PC_2, OUT_REG0,OUT_RESULT_ALU_1,OUT_MUX_MEM_TO_REG, NEW_MUX_SRC1_SEL, OUT_MUX_SRC1); --OUT_PC_2

MUX_ALU_SRC2 : MUX_5TO1 PORT MAP(OUT_REG_FILE2_1, OUT_IMM_GEN_1, OUT_REG4,OUT_RESULT_ALU_1,OUT_MUX_MEM_TO_REG, NEW_MUX_SRC2_SEL, OUT_MUX_SRC2);

MUX_OUT_MEM : MUX_2TO1 GENERIC MAP (64) PORT MAP(OUT_RESULT_ALU_2, DATA_OUT_MEM_DATA_1, MEM_TO_REG3, OUT_MUX_MEM_TO_REG );

RS1 <= INSTRUCTION_1(19 DOWNTO 15);
RS2 <= INSTRUCTION_1(24 DOWNTO 20);
RD <= INSTRUCTION_1(11 DOWNTO 7);

FORWARD_UNIT : ForwardingUnit PORT MAP (RS1_1, RS2_1, RD_2_EX_MEM, RD_3_MEM_WB,REG_WRITE2,REG_WRITE3,FORWARD_A,FORWARD_B,FA_FLAG,FB_FLAG);

Forward_on<=FA_FLAG OR FB_FLAG;

HAZARD_DETECTION : HazardDetectionUnit PORT MAP (RS1,RS2,RD_1,ADD_REG_WRITE_2,REG_WRITE3,MEM_READ1,Forward_on,CLK,EN_PC, EN_IF_ID, EN_ID_EX, MUX_SEL_BUBBLE);

EN_ISTR_MEM<=EN_IF_ID;

MUX_BUBBLE_OR_NOT : MUX_2TO1 GENERIC MAP (14) PORT MAP ("00000000000000",SIGNALS_CONTROL,MUX_SEL_BUBBLE,NEW_SIGNALS_CONTROL);

EN_FUNCT<=NEW_SIGNALS_CONTROL(13);
BRANCH <= NEW_SIGNALS_CONTROL(12);
MEM_READ <= NEW_SIGNALS_CONTROL(11); 
MEM_TO_REG <= NEW_SIGNALS_CONTROL(10); 
ALUop <= NEW_SIGNALS_CONTROL(9); 
MEM_WRITE <= NEW_SIGNALS_CONTROL(8); 
REG_WRITE <= NEW_SIGNALS_CONTROL(7);
MUX_TO_BRANCH <= NEW_SIGNALS_CONTROL(6);
ALU_src1 <= NEW_SIGNALS_CONTROL(5 DOWNTO 3);
ALU_src2 <= NEW_SIGNALS_CONTROL(2 DOWNTO 0);

MUX_FORWARD_CU_A : MUX_2TO1 GENERIC MAP (3) PORT MAP (ALU_src11, FORWARD_A, FA_FLAG, NEW_MUX_SRC1_SEL);

MUX_FORWARD_CU_B : MUX_2TO1 GENERIC MAP (3) PORT MAP (ALU_src21, FORWARD_B, FB_FLAG, NEW_MUX_SRC2_SEL);

MUX_BRANCH : MUX_2TO1 GENERIC MAP (1) PORT MAP(OUT_ZERO_ALU_1, (OTHERS=>'1'), MUX_TO_BRANCH2, OUT_MUX_BRANCH);

--(BIT(BRANCH3) AND BIT(OUT_MUX_BRANCH))

PROCESS(BRANCH2, OUT_MUX_BRANCH)

BEGIN

 IF(BRANCH2='1') THEN 

       IF(OUT_MUX_BRANCH="1") THEN SELECTOR_MUX_BRANCH_SEQ<='1';
		 
           ELSE SELECTOR_MUX_BRANCH_SEQ<='0';

			  END IF;
			  
   ELSE SELECTOR_MUX_BRANCH_SEQ<='0';

					 
  END IF;
  
END PROCESS;

MUX_BRANCH_SEQUENTIAL : MUX_2TO1 GENERIC MAP (64) PORT MAP(OUT_ADD_SEQUENTIAL, OUT_ADD_BRANCH_1, SELECTOR_MUX_BRANCH_SEQ, OUT_MUX_SEQ_BRANCH);

REG_0 : Register_N PORT MAP((OTHERS=>'0'),CLK, RST,'1', OUT_REG0);

REG_4 : Register_N PORT MAP(x"0000000000000004", CLK, RST,'1', OUT_REG4);




---------------------PIPE REGISTERS-------------


---------------------FIRST LEVEL---------------- 

PROCESS(CLK)
BEGIN
IF(CLK'EVENT AND CLK='1') THEN 
	IF(EN_IF_ID='1')THEN
	OUT_PC_1 <= OUT_MUX_PC; 
	ELSE 
	OUT_PC_1<=OUT_PC_1;
END IF;
END IF;
END PROCESS;


OUT_INSTR_FUNCT <= INSTRUCTION_1(14 DOWNTO 12);

--------------------SECOND LEVEL----------------

PROCESS(CLK)
BEGIN
IF(CLK'EVENT AND CLK='1') THEN 
	IF(EN_ID_EX='1') THEN 
	OPCODE_1<=INSTRUCTION_1(6 DOWNTO 0);
   ADD_REG_WRITE<=INSTRUCTION_1(11 DOWNTO 7);
   OUT_PC_2 <= OUT_PC_1; 
   OUT_REG_FILE1_1 <= OUT_REG_FILE1;
	OUT_REG_FILE2_1 <= OUT_REG_FILE2; 
	OUT_IMM_GEN_1 <= OUT_IMM_GEN; 
	OUT_INSTR_FUNCT_1 <= OUT_INSTR_FUNCT;
	RS1_1 <= RS1;
	RS2_1 <= RS2;
	RD_1 <=RD;
	ELSE 
	ADD_REG_WRITE<=ADD_REG_WRITE;
	OUT_PC_2 <= OUT_PC_2;  
	OUT_REG_FILE1_1 <= OUT_REG_FILE1_1;
	OUT_REG_FILE2_1 <= OUT_REG_FILE2_1; 
	OUT_IMM_GEN_1 <= OUT_IMM_GEN_1; 
	OUT_INSTR_FUNCT_1 <= OUT_INSTR_FUNCT_1;
	RS1_1 <= RS1_1;
	RS2_1 <= RS2_1;
	RD_1 <=RD_1;
	END IF;
END IF;
END PROCESS;

------------------------THIRD LEVEL--------------
 
PROCESS(CLK)
BEGIN
IF(CLK'EVENT AND CLK='1') THEN 
ADD_REG_WRITE_1<=ADD_REG_WRITE;
OUT_ADD_BRANCH_1 <= OUT_ADD_BRANCH;
OUT_ZERO_ALU_1 <= (OTHERS => OUT_ZERO_ALU);
OUT_RESULT_ALU_1 <= OUT_MUX_FUNCT_ALU; 
RD_2_EX_MEM <= RD_1;
END IF;
END PROCESS;



----------------------FOURTH LEVEL---------------


---REG WRITE, MEM TO REG
PROCESS(CLK)
BEGIN
IF(CLK'EVENT AND CLK='1') THEN 
ADD_REG_WRITE_2<=ADD_REG_WRITE_1;
DATA_OUT_MEM_DATA_1 <= DATA_OUT_MEM_DATA; 
OUT_RESULT_ALU_2 <= OUT_RESULT_ALU_1;
RD_3_MEM_WB <= RD_2_EX_MEM;
END IF;
END PROCESS;


--------------------------------------------PIPE CONTROLS-----------------------------------------


---------------------------------------FIRST LEVEL: ALL SIGNALS-----------------------------------
PROCESS(CLK)

BEGIN

IF(CLK'EVENT AND CLK='1') THEN 

BRANCH1 <= BRANCH; 
MEM_READ1 <= MEM_READ; 
MEM_WRITE1 <= MEM_WRITE; 
MEM_TO_REG1 <= MEM_TO_REG; 
ALUop1 <= ALUop; 
REG_WRITE1 <= REG_WRITE; 
MUX_TO_BRANCH1 <= MUX_TO_BRANCH; 
ALU_src11 <= ALU_src1; 
ALU_src21 <= ALU_src2;
EN_FUNCT1<=EN_FUNCT;

END IF;
END PROCESS;

--------------------------------------SECOND LEVEL ALL SIGNALS-------------------------------------
PROCESS(CLK)

BEGIN

IF(CLK'EVENT AND CLK='1') THEN 

BRANCH2 <= BRANCH1;  
MEM_TO_REG2 <= MEM_TO_REG1; 
REG_WRITE2 <= REG_WRITE1; 
MUX_TO_BRANCH2 <= MUX_TO_BRANCH1;

END IF;
END PROCESS;

READ_MEM_DATA<=MEM_READ1; 
WRITE_MEM_DATA<=MEM_WRITE1;
ADDRESS_MEM_DATA <= OUT_MUX_FUNCT_ALU;
DATA_TOWRITE_MEM_DATA <= OUT_REG_FILE2_1;

------------------------------------------THIRD LEVEL-----------------------------------
PROCESS(CLK)

BEGIN

IF(CLK'EVENT AND CLK='1') THEN 
 
MEM_TO_REG3 <= MEM_TO_REG2; 
REG_WRITE3 <= REG_WRITE2; 

END IF;
END PROCESS;

END ARCHITECTURE;


